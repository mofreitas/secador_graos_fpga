lpm_counterCONTADOR1_inst : lpm_counterCONTADOR1 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
