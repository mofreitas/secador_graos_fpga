library verilog;
use verilog.vl_types.all;
entity projeto3sd_vlg_vec_tst is
end projeto3sd_vlg_vec_tst;
